module rdy_valid_slave
#(parameter DW = 16)
